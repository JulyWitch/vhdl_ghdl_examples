LIBRARY ieee;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_ARITH.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY enc16x4 IS
    PORT (
        x : IN STD_LOGIC_VECTOR(15 DOWNTO 0);
        y : OUT STD_LOGIC_VECTOR(3 DOWNTO 0));

END enc16x4;

ARCHITECTURE rtl OF enc16x4 IS

BEGIN
    y <= "0000" WHEN (x = "0000000000000001") ELSE
        "0001" WHEN (x = "0000000000000010") ELSE
        "0010" WHEN (x = "0000000000000100") ELSE
        "0011" WHEN (x = "0000000000001000") ELSE
        "0100" WHEN (x = "0000000000010000") ELSE
        "0101" WHEN (x = "0000000000100000") ELSE
        "0110" WHEN (x = "0000000001000000") ELSE
        "0111" WHEN (x = "0000000010000000") ELSE
        "1000" WHEN (x = "0000000100000000") ELSE
        "1001" WHEN (x = "0000001000000000") ELSE
        "1010" WHEN (x = "0000010000000000") ELSE
        "1011" WHEN (x = "0000100000000000") ELSE
        "1100" WHEN (x = "0001000000000000") ELSE
        "1101" WHEN (x = "0010000000000000") ELSE
        "1110" WHEN (x = "0100000000000000") ELSE
        "1111" WHEN (x = "1000000000000000");

END ARCHITECTURE;